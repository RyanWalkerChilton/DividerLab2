library IEEE;
use IEEE.std_logic_1164.all;
--Additional standard or custom libraries go here if needed
package divider_const is
constant DIVIDEND_WIDTH:natural:=16;
constant DIVISOR_WIDTH:natural:=8;
end package body divider_const;